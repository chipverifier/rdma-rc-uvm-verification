package common_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
endpackage : common_pkg